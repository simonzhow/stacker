`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:10:13 06/02/2017 
// Design Name: 
// Module Name:    level 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module level(
	input clock,
	input [3:0] current_level,
	
	output [7:0] segment,
	output [3:0] an
	


    );


endmodule
